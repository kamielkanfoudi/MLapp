�csklearn.linear_model._logistic
LogisticRegression
q )�q}q(X   penaltyqX   l2qX   dualq�X   tolqG?6��C-X   CqG?�      X   fit_interceptq�X   intercept_scalingq	KX   class_weightq
NX   random_stateqNX   solverqX   lbfgsqX   max_iterqM�X   multi_classqX   multinomialqX   verboseqK X
   warm_startq�X   n_jobsqNX   l1_ratioqNX   n_features_in_qKX   classes_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   i8q���q Rq!(KX   <q"NNNJ����J����K tq#b�C               q$tq%bX   n_iter_q&hhK �q'h�q(Rq)(KK�q*hX   i4q+���q,Rq-(Kh"NNNJ����J����K tq.b�C�   q/tq0bX   coef_q1hhK �q2h�q3Rq4(KKK�q5hX   f8q6���q7Rq8(Kh"NNNJ����J����K tq9b�C�)��"w?�B.et��?�^R�%����d�i~;�?�c����t?a
g�h?�,%F�?�Tӵ��ֿ8��r��?�� ���^�`�d�;>�?�_v	��?�Жzߖο%�9/�m��v��	ʓ�?1l��Y�?{
[�ҽ?q:tq;bX
   intercept_q<hhK �q=h�q>Rq?(KK�q@h8�C��| �qAtqBbX   _sklearn_versionqCX   1.0.2qDub.